$date
  Mon Oct 10 22:27:07 2022
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module cont12b_lento_tb $end
$var reg 1 ! clk_t $end
$var reg 1 " rst_t $end
$var reg 1 # ena_t $end
$var reg 1 $ step_t $end
$var reg 1 % up_down_t $end
$var reg 12 & q_t[11:0] $end
$var reg 1 ' ena_o_t $end
$scope module int_cont $end
$var reg 1 ( clk_i $end
$var reg 1 ) rst_i $end
$var reg 1 * ena_i $end
$var reg 1 + step_i $end
$var reg 1 , up_down $end
$var reg 12 - q_o[11:0] $end
$var reg 1 . ena_o $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
0!
1"
1#
0$
0%
bUUUUUUUUUUUU &
U'
0(
1)
1*
0+
0,
bUUUUUUUUUUUU -
U.
#10000000
1!
b000000000000 &
0'
1(
b000000000000 -
0.
#20000000
0!
0(
#30000000
1!
1(
#40000000
0!
0(
#50000000
1!
0"
1(
0)
#60000000
0!
0(
#70000000
1!
b000000000001 &
1'
1(
b000000000001 -
1.
#80000000
0!
0(
#90000000
1!
0'
1(
0.
#100000000
0!
0(
#110000000
1!
b000000000010 &
1'
1(
b000000000010 -
1.
#120000000
0!
0(
#130000000
1!
0'
1(
0.
#140000000
0!
0(
#150000000
1!
b000000000011 &
1'
1(
b000000000011 -
1.
#160000000
0!
0(
#170000000
1!
0'
1(
0.
#180000000
0!
0(
#190000000
1!
b000000000100 &
1'
1(
b000000000100 -
1.
#200000000
0!
0(
#210000000
1!
0'
1(
0.
#220000000
0!
0(
#230000000
1!
b000000000101 &
1'
1(
b000000000101 -
1.
#240000000
0!
0(
#250000000
1!
0'
1(
0.
#260000000
0!
0(
#270000000
1!
b000000000110 &
1'
1(
b000000000110 -
1.
#280000000
0!
0(
#290000000
1!
0'
1(
0.
#300000000
0!
0(
#310000000
1!
b000000000111 &
1'
1(
b000000000111 -
1.
#320000000
0!
0(
#330000000
1!
0'
1(
0.
#340000000
0!
0(
#350000000
1!
b000000001000 &
1'
1(
b000000001000 -
1.
#360000000
0!
0(
#370000000
1!
0'
1(
0.
#380000000
0!
0(
#390000000
1!
b000000001001 &
1'
1(
b000000001001 -
1.
#400000000
0!
0(
#410000000
1!
0'
1(
0.
#420000000
0!
0(
#430000000
1!
b000000001010 &
1'
1(
b000000001010 -
1.
#440000000
0!
0(
#450000000
1!
0'
1(
0.
#460000000
0!
0(
#470000000
1!
b000000001011 &
1'
1(
b000000001011 -
1.
#480000000
0!
0(
#490000000
1!
0'
1(
0.
#500000000
0!
1$
0(
1+
#510000000
1!
b000000001101 &
1'
1(
b000000001101 -
1.
#520000000
0!
0(
#530000000
1!
0'
1(
0.
#540000000
0!
0(
#550000000
1!
b000000001111 &
1'
1(
b000000001111 -
1.
#560000000
0!
0(
#570000000
1!
0'
1(
0.
#580000000
0!
0(
#590000000
1!
b000000010001 &
1'
1(
b000000010001 -
1.
#600000000
0!
0(
#610000000
1!
0'
1(
0.
#620000000
0!
0#
0(
0*
#630000000
1!
1(
#640000000
0!
0(
#650000000
1!
1(
#660000000
0!
0(
#670000000
1!
1(
#680000000
0!
0(
#690000000
1!
1(
#700000000
0!
0(
#710000000
1!
1(
#720000000
0!
0(
#730000000
1!
1(
#740000000
0!
0(
#750000000
1!
1(
#760000000
0!
0(
#770000000
1!
1(
#780000000
0!
0(
#790000000
1!
1(
#800000000
0!
1#
0(
1*
#810000000
1!
b000000010011 &
1'
1(
b000000010011 -
1.
#820000000
0!
0(
#830000000
1!
0'
1(
0.
#840000000
0!
0(
#850000000
1!
b000000010101 &
1'
1(
b000000010101 -
1.
#860000000
0!
0(
#870000000
1!
0'
1(
0.
#880000000
0!
0(
#890000000
1!
b000000010111 &
1'
1(
b000000010111 -
1.
#900000000
0!
0(
#910000000
1!
0'
1(
0.
#920000000
0!
0(
#930000000
1!
b000000011001 &
1'
1(
b000000011001 -
1.
#940000000
0!
0(
#950000000
1!
0'
1(
0.
#960000000
0!
0(
#970000000
1!
b000000011011 &
1'
1(
b000000011011 -
1.
#980000000
0!
0(
#990000000
1!
0'
1(
0.
#1000000000
0!
0$
0(
0+
#1010000000
1!
b000000011100 &
1'
1(
b000000011100 -
1.
#1020000000
0!
0(
#1030000000
1!
0'
1(
0.
#1040000000
0!
0(
#1050000000
1!
b000000011101 &
1'
1(
b000000011101 -
1.
#1060000000
0!
0(
#1070000000
1!
0'
1(
0.
#1080000000
0!
0(
#1090000000
1!
b000000011110 &
1'
1(
b000000011110 -
1.
#1100000000
0!
0(
#1110000000
1!
0'
1(
0.
#1120000000
0!
0(
#1130000000
1!
b000000011111 &
1'
1(
b000000011111 -
1.
#1140000000
0!
0(
#1150000000
1!
0'
1(
0.
#1160000000
0!
0(
#1170000000
1!
b000000100000 &
1'
1(
b000000100000 -
1.
#1180000000
0!
0(
#1190000000
1!
0'
1(
0.
#1200000000
0!
0(
#1210000000
1!
b000000100001 &
1'
1(
b000000100001 -
1.
#1220000000
0!
0(
#1230000000
1!
0'
1(
0.
#1240000000
0!
0(
#1250000000
1!
b000000100010 &
1'
1(
b000000100010 -
1.
#1260000000
0!
0(
#1270000000
1!
0'
1(
0.
#1280000000
0!
0(
#1290000000
1!
b000000100011 &
1'
1(
b000000100011 -
1.
#1300000000
0!
1%
0(
1,
#1310000000
1!
0'
1(
0.
#1320000000
0!
0(
#1330000000
1!
b000000100010 &
1'
1(
b000000100010 -
1.
#1340000000
0!
0(
#1350000000
1!
0'
1(
0.
#1360000000
0!
0(
#1370000000
1!
b000000100001 &
1'
1(
b000000100001 -
1.
#1380000000
0!
0(
#1390000000
1!
0'
1(
0.
#1400000000
0!
0(
#1410000000
1!
b000000100000 &
1'
1(
b000000100000 -
1.
#1420000000
0!
0(
#1430000000
1!
0'
1(
0.
#1440000000
0!
0(
#1450000000
1!
b000000011111 &
1'
1(
b000000011111 -
1.
#1460000000
0!
0(
#1470000000
1!
0'
1(
0.
#1480000000
0!
0(
#1490000000
1!
b000000011110 &
1'
1(
b000000011110 -
1.
#1500000000
0!
1$
0(
1+
#1510000000
1!
0'
1(
0.
#1520000000
0!
0(
#1530000000
1!
b000000011100 &
1'
1(
b000000011100 -
1.
#1540000000
0!
0(
#1550000000
1!
0'
1(
0.
#1560000000
0!
0(
#1570000000
1!
b000000011010 &
1'
1(
b000000011010 -
1.
#1580000000
0!
0(
#1590000000
1!
0'
1(
0.
#1600000000
0!
0(
#1610000000
1!
b000000011000 &
1'
1(
b000000011000 -
1.
#1620000000
0!
0(
#1630000000
1!
0'
1(
0.
#1640000000
0!
0(
#1650000000
1!
b000000010110 &
1'
1(
b000000010110 -
1.
#1660000000
0!
0(
#1670000000
1!
0'
1(
0.
#1680000000
0!
0(
#1690000000
1!
b000000010100 &
1'
1(
b000000010100 -
1.
#1700000000
0!
0(
#1710000000
1!
0'
1(
0.
#1720000000
0!
0(
#1730000000
1!
b000000010010 &
1'
1(
b000000010010 -
1.
#1740000000
0!
0(
#1750000000
1!
0'
1(
0.
#1760000000
0!
0(
#1770000000
1!
b000000010000 &
1'
1(
b000000010000 -
1.
#1780000000
0!
0(
#1790000000
1!
0'
1(
0.
#1800000000
0!
0(
#1810000000
1!
b000000001110 &
1'
1(
b000000001110 -
1.
#1820000000
0!
0(
#1830000000
1!
0'
1(
0.
#1840000000
0!
0(
#1850000000
1!
b000000001100 &
1'
1(
b000000001100 -
1.
#1860000000
0!
0(
#1870000000
1!
0'
1(
0.
#1880000000
0!
0(
#1890000000
1!
b000000001010 &
1'
1(
b000000001010 -
1.
#1900000000
0!
0(
#1910000000
1!
0'
1(
0.
#1920000000
0!
0(
#1930000000
1!
b000000001000 &
1'
1(
b000000001000 -
1.
#1940000000
0!
0(
#1950000000
1!
0'
1(
0.
#1960000000
0!
0(
#1970000000
1!
b000000000110 &
1'
1(
b000000000110 -
1.
#1980000000
0!
0(
#1990000000
1!
0'
1(
0.
#2000000000
0!
0(
